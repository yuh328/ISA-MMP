3&u��K9�D{n���rf��5uڴ��#�+q�0r�%}K��-����Wt�~��/��$[+v��+���Nk�#�+�u(�l�4����ơ��8��iL�od	�yY��ڊ	��5IAܕp���)/�"}�cHW@)蚼���oL�$6U&�=��p� �����,h&�kӋ�DR�h��ҞX~[�\��[ɧ�>'���,]�!d���#����"\ZH.=%.��i�c��<f�z�o��Z����		UL/�sB��%��$�V��X��������1W�T�578;�L�;�2�f����� ��w=�Z�\���G���d�N�]/Z��M�C��� �e�p����+G<���b��Y�����KY���|���s)��i������oVe�?1�t����P.����9�sr��ZKȋV�� Έ�Â���6��O7��^?A����B��P��`#��E2M�AY�M<�eq����S)pE�3xl�|���7&Ĺ��\�ܹR<XZC���W��%�Ƌ!^�LI�a�AS�9�j{dQ�KYo��f�����!���pj-V���;�V�q��alx��������n�#�ABu�r�+d��T��0k�qs��t�/