^2b������:���H��D9�R9c�AU|V=��<}��36|G���� ���{��o�߫�D�^���o}֭�̖u����k!Լ
z/��̖�~^N���d/R԰��m22nܜ͛�Cx���_|c`�ba��	�D�����B(��k��D�2�dz}ּ۪��}^��I. �2����=���e���~i�sG*�i������α�J֎}�g�eU1R����w5P��[��a�[.����=�1���r�����d��:?θ�]kÆF������/�~G��#���y����;���Z��]3������s�� �q���"����Wv!��و�T���"�����T�������PP�f��CNUl�O�RMDv�:�i�������<��5�@J��8��*\����jj@`�᳢�@�a��;	��og�1��